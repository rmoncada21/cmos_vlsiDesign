// Created Sun Dec  1 11:52:56 2024

module flipflop_1bit ();

  always begin
	test
  end
endmodule
