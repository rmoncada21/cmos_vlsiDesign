* libro_models.sp
**---------------------------------------------------------
* Modelos NMOS y PMOS
**---------------------------------------------------------
.model NMOS NMOS (LEVEL=1 VTO=0.7 KP=120u LAMBDA=0.02)
.model PMOS PMOS (LEVEL=1 VTO=-0.7 KP=50u LAMBDA=0.02)
